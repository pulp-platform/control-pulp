/*
 * pulp_soc_defines.sv
 *
 * Copyright (C) 2013-2018 ETH Zurich, University of Bologna.
 *
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 */

`ifndef PULP_SOC_DEFINES_SV
`define PULP_SOC_DEFINES_SV

// define if the 0x0000_0000 to 0x0040_0000 is the alias of the current cluster
// address space (eg cluster 0 is from 0x1000_0000 to 0x1040_0000)
`define CLUSTER_ALIAS
// the same for fabric controller
`define FC_ALIAS

// To use new icache use this define
//`define MP_ICACHE
//`define SP_ICACHE
`define PRIVATE_ICACHE
`define HIERARCHY_ICACHE_32BIT

// To use The L2 Multibank Feature, please decomment this define
`define USE_L2_MULTIBANK
`define NB_L2_CHANNELS 4


// JTAG
// Part Number
//   0001/fffe PULPissimo
//   0002/fffd PULP
//   cafe/3501 ControlPULP

// LSB                       [0]:     1'h1
// PULP Platform Manufacturer[11:1]:  11'h6d9
// Part Number               [27:12]: 16'hcafe
// Version                   [31:28]: 4'h5
`define DMI_JTAG_IDCODE 32'h5cafedb3

// LSB                       [0]:     1'h1
// PULP Platform Manufacturer[11:1]:  11'h6d9
// Part Number               [27:12]: 16'hcaff
// Version                   [31:28]: 4'h5
`define PULP_JTAG_IDCODE 32'h53501db3


// FPU
`define FPU_CLUSTER

// Debugging
// Trace CV32E40P core execution
// `define CV32E40P_TRACE_EXECUTION
// Trace CV32E40P offload interface
// `define CV32E40P_APU_TRACE
// Compare the output of the instruction CACHE with the slm files generated by the compiler
//`define DEBUG_FETCH_INTERFACE
// Log soc, peripheral and cluster clock frequencies
//`define DEBUG_CLK_RST_GEN
// Log uart output
`define LOG_UART_SIM
// Log sim stdout to files
//`define LOG_SIM_STDOUT


// If you want to place the DEMUX peripherals (EU, MCHAN) rigth before the Test and set region.
// This will steal 16KB from the 1MB TCDM reegion.
// EU is mapped           from 0x10100000 - 0x400
// MCHAN regs are mapped  from 0x10100000 - 0x800
//`define DEM_PER_BEFORE_TCDM_TS

// Enables memory mapped register and counters to extract statistic on instruction cache
`define FEATURE_ICACHE_STAT

// Parameters
`define NB_CLUSTERS      1
`define NB_CORES         8
`define DMA_QUEUE_DEPTH  8
`define TWD_QUEUE_DEPTH  4
`define NB_DMAS          4
`define NB_OUTSND_BURSTS 16
`define NB_MPERIPHS      1
`define NB_SPERIPHS      10
`define GPIO_NUM         64

// Width of byte enable for a given data width
`define EVAL_BE_WIDTH(DATAWIDTH) (DATAWIDTH/8)

// Helpers
`define LOG2(VALUE) ((VALUE) < ( 1 ) ? 0 : (VALUE) < ( 2 ) ? 1 : (VALUE) < ( 4 ) ? 2 : (VALUE)< (8) ? 3:(VALUE) < ( 16 )  ? 4 : (VALUE) < ( 32 )  ? 5 : (VALUE) < ( 64 )  ? 6 : (VALUE) < ( 128 ) ? 7 : (VALUE) < ( 256 ) ? 8 : (VALUE) < ( 512 ) ? 9 : 10)

`endif
